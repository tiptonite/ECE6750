library IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.NUMERIC_STD.all;
package bus_multiplier_pkg is
        type bus_array is array(0 to 127 ) of unsigned(7 downto 0);
end package;